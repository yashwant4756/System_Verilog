module array_problem;
  import "DPI-C" context function void arr();
  initial run();
 task run();
     arr();
   endtask
endmodule
